library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package Common is

	type Q_array is array(0 to 15) of std_logic_vector(11 downto 0);

end Common;

package body Common is
   -- subprogram bodies here
end Common;